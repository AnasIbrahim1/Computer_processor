/*******************************************************************
*
* Module: ProcessorMain.v
* Project: Processor
* Authors: Anas A. Ibrahim - anas2@aucegypt.edu, Ibrahim Gohar - 
abdelmaksou@aucegypt.edu

* Description: main processor circuit, where all the modules are combined
*
* Change history: 06/11/2022 - Added from Lab 6
                  06/11/2022 - Additional gates/muxes/modules were added to support all
                  instruction
                  13/11/2022 - Creation Date
			21/11/2022 - Updated out and mem_out to avoid Don't Care
*
**********************************************************************/
module SingleMem(
    input is_inst,
    input MemRead, 
    input MemWrite,
    input [2 : 0] funct3,
    input [8  : 0] addr, 
    input [31 : 0] in, 
    output reg[31 : 0] out,
    output reg[31 : 0] mem_out
);

    reg[7 : 0] mem[511 : 0];
    wire[8 : 0] new_addr;
    assign new_addr = { addr[7 : 0], is_inst };
    // data are even and instructions are odd
     always @(*) begin
        if (is_inst) begin
            out <= {mem[new_addr + 6], mem[new_addr + 4], mem[new_addr + 2], mem[new_addr + 0]};
            mem_out <= mem_out;
        end else begin
            if (MemWrite) begin 
                if (funct3 == `LS_FUNCT3_B) 
                    mem[new_addr] <= in[7 : 0];
                else if (funct3 == `LS_FUNCT3_H) begin
                    mem[new_addr] <= in[7 : 0];
                    mem[new_addr + 2] <= in[15 : 8];                
                end else begin
                    mem[new_addr] <= in[7 : 0];
                    mem[new_addr + 2] <= in[15 : 8];                
                    mem[new_addr + 4] <= in[23 : 16];
                    mem[new_addr + 6] <= in[31 : 24];                
                end
                mem_out <= mem_out;
            end 
            else if (MemRead) begin
                if (funct3 == `LS_FUNCT3_B) 
                    mem_out <= { { 24 { mem[new_addr][7] } }, mem[new_addr] };
                else if (funct3 == `LS_FUNCT3_H) 
                    mem_out <= { { 16 { mem[new_addr + 2][7] } }, mem[new_addr + 2], mem[new_addr] };
                else if (funct3 == `LS_FUNCT3_BU) 
                    mem_out <= { 24'b0 , mem[new_addr] };
                else if (funct3 == `LS_FUNCT3_HU) 
                    mem_out <= { 16'b0 , mem[new_addr + 2], mem[new_addr] };
                else 
                    mem_out <= { mem[new_addr + 6], mem[new_addr + 4], mem[new_addr + 2], mem[new_addr] };
            end
            out <= out;
        end
    end
    
    parameter nop = 32'b0000000_00000_00000_000_00000_0110011;
    initial begin
    // memory data
        {mem[6], mem[4], mem[2], mem[0]} = 32'd17;
        {mem[14], mem[12], mem[10], mem[8]} = 32'd9;
        {mem[22], mem[20], mem[18], mem[16]} = 32'd25;

           // inst data

// With NOPS
         
//            {mem[7], mem[5], mem[3], mem[1]}         = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[15], mem[13], mem[11], mem[9]}      = 32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0)
//            {mem[23], mem[21], mem[19], mem[17]}      = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[31], mem[29], mem[27], mem[25]}      = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[39], mem[37], mem[35], mem[33]}      = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[47], mem[45], mem[43], mem[41]}      = 32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)
//            {mem[55], mem[53], mem[51], mem[49]}       = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[63], mem[61], mem[59], mem[57]}      = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[71], mem[69], mem[67], mem[65]}      = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[79], mem[77], mem[75], mem[73]}      = 32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0)
//            {mem[87], mem[85], mem[83], mem[81]}     = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[95], mem[93], mem[91], mem[89]}     = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[103], mem[101], mem[99], mem[97]}  = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[111], mem[109], mem[107], mem[105]} = 32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2
//            {mem[119], mem[117], mem[115], mem[113]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[127], mem[125], mem[123], mem[121]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[135], mem[133], mem[131], mem[129]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[143], mem[141], mem[139], mem[137]} = 32'b0_000001_00011_00100_000_0000_0_1100011; //beq x4, x3, 16
//            {mem[151], mem[149], mem[147], mem[145]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[159], mem[157], mem[155], mem[153]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[167], mem[165], mem[163], mem[161]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[175], mem[173], mem[171], mem[169]} = 32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2
//            {mem[183], mem[181], mem[179], mem[177]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[191], mem[189], mem[187], mem[185]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[199], mem[197], mem[195], mem[193]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[207], mem[205], mem[203], mem[201]}= 32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2
//            {mem[215], mem[213], mem[211], mem[209]}= 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[223], mem[221], mem[219], mem[217]}= 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[231], mem[229], mem[227], mem[225]}= 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0  
//            {mem[239], mem[237], mem[235], mem[233]}= 32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)
//            {mem[247], mem[245], mem[243], mem[241]}= 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[255], mem[253], mem[251], mem[249]}= 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[263], mem[261], mem[259], mem[257]}= 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[271], mem[269], mem[267], mem[265]}= 32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
//            {mem[279], mem[277], mem[275], mem[273]}= 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[287], mem[285], mem[283], mem[281]}= 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[295], mem[293], mem[291], mem[289]}= 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[303], mem[301], mem[299], mem[297]}= 32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1
//            {mem[311], mem[309], mem[307], mem[305]}= 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[319], mem[317], mem[315], mem[313]}= 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[327], mem[325], mem[323], mem[321]}= 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[335], mem[333], mem[331], mem[329]}= 32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2
//            {mem[343], mem[341], mem[339], mem[337]}= 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[351], mem[349], mem[347], mem[345]}= 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[359], mem[357], mem[355], mem[353]}= 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[367], mem[365], mem[363], mem[361]} = 32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2
//            {mem[375], mem[373], mem[371], mem[369]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[383], mem[381], mem[379], mem[377]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[391], mem[389], mem[387], mem[385]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[399], mem[397], mem[395], mem[393]} = 32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1
//            {mem[407], mem[405], mem[403], mem[401]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[415], mem[413], mem[411], mem[409]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
//            {mem[423], mem[421], mem[419], mem[417]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0

           
// NO NOPS
             
           /*
           {mem[7], mem[5], mem[3], mem[1]}          = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
           {mem[15], mem[13], mem[11], mem[9]}       = 32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0)
           {mem[23], mem[21], mem[19], mem[17]}      = 32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)
           {mem[31], mem[29], mem[27], mem[25]}      = 32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0)
           {mem[39], mem[37], mem[35], mem[33]}      = 32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2
           {mem[47], mem[45], mem[43], mem[41]}      = 32'h00320463; //beq x4, x3, 8                                 
           {mem[55], mem[53], mem[51], mem[49]}      = 32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2    
           {mem[63], mem[61], mem[59], mem[57]}      = 32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2    
           {mem[71], mem[69], mem[67], mem[65]}      = 32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)   
           {mem[79], mem[77], mem[75], mem[73]}      = 32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)   
           {mem[87], mem[85], mem[83], mem[81]}      = 32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1 
           {mem[95], mem[93], mem[91], mem[89]}      = 32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2 
           {mem[103], mem[101], mem[99], mem[97]}    = 32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2 
           {mem[111], mem[109], mem[107], mem[105]}  = 32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1 

		*/

    end    
endmodule
